module pacmanrom ( input [6:0]	addr,
				  output [12:0]	data
					 );

	parameter ADDR_WIDTH = 7;
	parameter DATA_WIDTH =  13;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	   //code x00
	   13'b0000111110000,
	   13'b0011111111100,
	   13'b0111111111110,
	   13'b0111111111110,
	   13'b1111111111111,
	   13'b1111111111111,
	   13'b1111111111111,
	   13'b1111111111111,
	   13'b1111111111111,
	   13'b0111111111110,
	   13'b0111111111110,
	   13'b0011111111100,
	   13'b0000111110000,
	   
	   //code x01
	   13'b0000000000000,
	   13'b0011000001100,
	   13'b0111000001110,
	   13'b0111100011110,
	   13'b1111100011111,
	   13'b1111100011111,
	   13'b1111110111111,
	   13'b1111110111111,
	   13'b1111110111111,
	   13'b0111111111110,
	   13'b0111111111110,
	   13'b0011111111100,
	   13'b0000111110000,
	   
	   //code x02
	   13'b0000000000000,
	   13'b0000000000000,
	   13'b0000000000000,
	   13'b0000000000000,
	   13'b1100000000011,
	   13'b1110000000111,
	   13'b1111000001111,
	   13'b1111100011111,
	   13'b1111110111111,
	   13'b0111111111110,
	   13'b0111111111110,
	   13'b0011111111100,
	   13'b0000111110000,
	   
	   //code x03
	   13'b0000111110000,
	   13'b0011111111100,
	   13'b0111111111110,
	   13'b0111111111110,
	   13'b1111111111000,
	   13'b1111110000000,
	   13'b1111000000000,
	   13'b1111110000000,
	   13'b1111111111000,
	   13'b0111111111110,
	   13'b0111111111110,
       13'b0011111111100,
       13'b0000111110000,
       
       
       //code x04
       13'b0000111110000,
       13'b0011111110000,
       13'b0111111100000,
       13'b0111111000000,
       13'b1111110000000,
       13'b1111100000000,
       13'b1111000000000,
       13'b1111100000000,
       13'b1111110000000,
       13'b0111111000000,
       13'b0111111100000,
       13'b0011111110000,
       13'b0000111110000,
       
       //code x05
       13'b0000111110000,
       13'b0011111111100,
       13'b0111111111110,
       13'b0111111111110,
       13'b1111110111111,
       13'b1111110111111,
       13'b1111110111111,
       13'b1111100011111,
       13'b1111100011111,
       13'b0111100011110,
       13'b0111000001110,
       13'b0011000001100,
       13'b0000000000000,
       
       //code x06
       13'b0000111110000,
       13'b0011111111100,
       13'b0111111111110,
       13'b0111111111110,
       13'b1111110111111,
       13'b1111100011111,
       13'b1111000001111,
       13'b1110000000111,
       13'b1100000000011,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       
       //code x07
       13'b0000111110000,
       13'b0011111111100,
       13'b0111111111110,
       13'b0111111111110,
       13'b0001111111111,
       13'b0000001111111,
       13'b0000000001111,
       13'b0000001111111,
       13'b0001111111111,
       13'b0111111111110,
       13'b0111111111110,
       13'b0011111111100,
       13'b0000111110000,
       
       //code x08
       13'b0000111110000,
       13'b0000111111100,
       13'b0000011111110,
       13'b0000001111110,
       13'b0000000111111,
       13'b0000000011111,
       13'b0000000001111,
       13'b0000000011111,
       13'b0000000111111,
       13'b0000001111110,
       13'b0000011111110,
       13'b0000111111100,
       13'b0000111110000,
       
       //xx
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000,
       13'b0000000000000 
      };

	assign data = ROM[addr];

endmodule  
