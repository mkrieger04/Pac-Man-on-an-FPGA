module ghostfont ( input [4:0]	addr,
				  output [27:0]	data
					 );

	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH =  28;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	   //code x01
      28'b0000000000111111110000000000,
      28'b0000001111111111111111000000,
      28'b0000111111111111111111110000,
      28'b0011110101111111110101111100,
      28'b0011010101011111010101011100,
      28'b0011011010011111011010011100,
      28'b1111011010011111011010011111,           
      28'b1111110101111111110101111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111001111110000111111001111,
      28'b1100000011110000111100000011,
      //code 2
      28'b0000000000111111110000000000,
      28'b0000001111111111111111000000,
      28'b0000111111111111111111110000,
      28'b0011110101111111110101111100,
      28'b0011010101011111010101011100,
      28'b0011011010011111011010011100,
      28'b1111011010011111011010011111,           
      28'b1111110101111111110101111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111111111111111111111111111,
      28'b1111111100111111110011111111,
      28'b1111110000001111000000111111,
      
      //yuck
      28'b0000000000000000000000000000,
      28'b0000000000000000000000000000,
      28'b0000000000000000000000000000,
      28'b0000000000000000000000000000
      
      };

	assign data = ROM[addr];

endmodule  
